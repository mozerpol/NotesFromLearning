     a_in <= '0';
     b_in <= '0';
     wait for 1 us;
