module tff(
   input wire clk,
   input wire t,
   output wire q
);
endmodule
