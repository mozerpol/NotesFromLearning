library ieee;
   use ieee.std_logic_1164.all;


 package my_design_pkg is


   constant C_DATA_WIDTH  : integer := 5;


 end;


 package body my_design_pkg is


 end package body;
