module dff(
   input wire clk,
   input wire d,
   output wire q
);
endmodule
