module simpleRAM #(
   parameter wordSize = 8,
   parameter addressSize = 32
)(
   input wire clk,
   input wire we,
   input wire re,
   inout wire data
);
endmodule
