module jkff(
   input wire clk,
   input wire j,
   input wire k,
   output wire q
);
endmodule
