     a_in <= 'Z';
     b_in <= 'Z';
     wait for 1 us;
