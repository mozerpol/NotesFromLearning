module srff(
   input wire clk,
   input wire s,
   input wire r,
   output wire q
);



endmodule
