library ieee;
  use ieee.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;
  
 package simplegate_pkg is
    constant C_TEST : std_logic_vector(1 downto 0) := "11";
 end;
 
 package body simplegate_pkg is
 
 end package body;
