module counter #(
   parameter N = 10
)(
   input wire clk,
   input wire rst,
   input wire ce,
   output wire ov
);
   
   

endmodule
