     a_in <= '1';
     b_in <= '1';
     wait for 1 us;
