library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.math_real.all;
  
 package and_gate_pkg is
    constant C_TEST : std_logic_vector(1 downto 0) := "11";
 end;
 
 package body and_gate_pkg is
 
 end package body;
