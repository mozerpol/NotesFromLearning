module uart_tx
	#(parameter BAUD = 9600)
	(
	input clk,
	input rst,
	input [7:0] data,
	output tx
);


endmodule
