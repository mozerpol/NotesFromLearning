library ieee;
  use ieee.std_logic_1164.all;

entity and_area is port (
    in1      : in    std_logic;
    in2      : in    std_logic;
    out1_and : out   std_logic
  );
end entity and_area;

architecture rtl of and_area is

begin

  and_process : process is
  begin

  end process and_process;

end architecture rtl;
