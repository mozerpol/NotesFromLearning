library ieee;
   use ieee.std_logic_1164.all;


package all_gates_pkg is
   constant C_TEST : std_logic_vector(1 downto 0) := "11";
end;


package body all_gates_pkg is


end package body;
