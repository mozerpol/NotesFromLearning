module uart_rx #(
   parameter F = 8000000,
   parameter BAUD = 115200
) (
   input wire rx
);
endmodule
